----------------------------------------------------------------------------------------------------
-- Copyright (c) 2023 Marcus Geelnard
--
-- This software is provided 'as-is', without any express or implied warranty. In no event will the
-- authors be held liable for any damages arising from the use of this software.
--
-- Permission is granted to anyone to use this software for any purpose, including commercial
-- applications, and to alter it and redistribute it freely, subject to the following restrictions:
--
--  1. The origin of this software must not be misrepresented; you must not claim that you wrote
--     the original software. If you use this software in a product, an acknowledgment in the
--     product documentation would be appreciated but is not required.
--
--  2. Altered source versions must be plainly marked as such, and must not be misrepresented as
--     being the original software.
--
--  3. This notice may not be removed or altered from any source distribution.
----------------------------------------------------------------------------------------------------

----------------------------------------------------------------------------------------------------
-- This implements CRC-32C (Castagnoli), polynomial 0x1edc6f41.
--
-- CRC polynomial coefficients: x^32 + x^28 + x^27 + x^26 + x^25 + x^23 + x^22 + x^20 + x^19 +
--                              x^18 + x^14 + x^13 + x^11 + x^10 + x^9 + x^8 + x^6 + 1
--
-- Combinatorial logic generated by: https://bues.ch/h/crcgen
----------------------------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use work.types.all;
use work.config.all;

entity crc32c is
  port (
    i_crc: in std_logic_vector(31 downto 0);
    i_data: in std_logic_vector(31 downto 0);
    i_packed_mode : in T_PACKED_MODE;
    o_result: out std_logic_vector(31 downto 0)
  );
end crc32c;

architecture rtl of crc32c is
  signal s_result8 : std_logic_vector(31 downto 0);
  signal s_result16 : std_logic_vector(31 downto 0);
  signal s_result32 : std_logic_vector(31 downto 0);
begin
  -- 8 bits per clock (only bits 7 downto 0 are used from i_data).
  s_result8(0) <= (i_crc(0) xor i_crc(1) xor i_crc(2) xor i_crc(3) xor i_crc(4) xor i_crc(8) xor i_data(0) xor i_data(1) xor i_data(2) xor i_data(3) xor i_data(4));
  s_result8(1) <= (i_crc(0) xor i_crc(1) xor i_crc(2) xor i_crc(3) xor i_crc(4) xor i_crc(5) xor i_crc(9) xor i_data(0) xor i_data(1) xor i_data(2) xor i_data(3) xor i_data(4) xor i_data(5));
  s_result8(2) <= (i_crc(1) xor i_crc(2) xor i_crc(3) xor i_crc(4) xor i_crc(5) xor i_crc(6) xor i_crc(10) xor i_data(1) xor i_data(2) xor i_data(3) xor i_data(4) xor i_data(5) xor i_data(6));
  s_result8(3) <= (i_crc(2) xor i_crc(3) xor i_crc(4) xor i_crc(5) xor i_crc(6) xor i_crc(7) xor i_crc(11) xor i_data(2) xor i_data(3) xor i_data(4) xor i_data(5) xor i_data(6) xor i_data(7));
  s_result8(4) <= (i_crc(1) xor i_crc(2) xor i_crc(5) xor i_crc(6) xor i_crc(7) xor i_crc(12) xor i_data(1) xor i_data(2) xor i_data(5) xor i_data(6) xor i_data(7));
  s_result8(5) <= (i_crc(1) xor i_crc(4) xor i_crc(6) xor i_crc(7) xor i_crc(13) xor i_data(1) xor i_data(4) xor i_data(6) xor i_data(7));
  s_result8(6) <= (i_crc(1) xor i_crc(3) xor i_crc(4) xor i_crc(5) xor i_crc(7) xor i_crc(14) xor i_data(1) xor i_data(3) xor i_data(4) xor i_data(5) xor i_data(7));
  s_result8(7) <= (i_crc(1) xor i_crc(3) xor i_crc(5) xor i_crc(6) xor i_crc(15) xor i_data(1) xor i_data(3) xor i_data(5) xor i_data(6));
  s_result8(8) <= (i_crc(0) xor i_crc(2) xor i_crc(4) xor i_crc(6) xor i_crc(7) xor i_crc(16) xor i_data(0) xor i_data(2) xor i_data(4) xor i_data(6) xor i_data(7));
  s_result8(9) <= (i_crc(0) xor i_crc(2) xor i_crc(4) xor i_crc(5) xor i_crc(7) xor i_crc(17) xor i_data(0) xor i_data(2) xor i_data(4) xor i_data(5) xor i_data(7));
  s_result8(10) <= (i_crc(2) xor i_crc(4) xor i_crc(5) xor i_crc(6) xor i_crc(18) xor i_data(2) xor i_data(4) xor i_data(5) xor i_data(6));
  s_result8(11) <= (i_crc(3) xor i_crc(5) xor i_crc(6) xor i_crc(7) xor i_crc(19) xor i_data(3) xor i_data(5) xor i_data(6) xor i_data(7));
  s_result8(12) <= (i_crc(1) xor i_crc(2) xor i_crc(3) xor i_crc(6) xor i_crc(7) xor i_crc(20) xor i_data(1) xor i_data(2) xor i_data(3) xor i_data(6) xor i_data(7));
  s_result8(13) <= (i_crc(1) xor i_crc(7) xor i_crc(21) xor i_data(1) xor i_data(7));
  s_result8(14) <= (i_crc(1) xor i_crc(3) xor i_crc(4) xor i_crc(22) xor i_data(1) xor i_data(3) xor i_data(4));
  s_result8(15) <= (i_crc(0) xor i_crc(2) xor i_crc(4) xor i_crc(5) xor i_crc(23) xor i_data(0) xor i_data(2) xor i_data(4) xor i_data(5));
  s_result8(16) <= (i_crc(0) xor i_crc(1) xor i_crc(3) xor i_crc(5) xor i_crc(6) xor i_crc(24) xor i_data(0) xor i_data(1) xor i_data(3) xor i_data(5) xor i_data(6));
  s_result8(17) <= (i_crc(0) xor i_crc(1) xor i_crc(2) xor i_crc(4) xor i_crc(6) xor i_crc(7) xor i_crc(25) xor i_data(0) xor i_data(1) xor i_data(2) xor i_data(4) xor i_data(6) xor i_data(7));
  s_result8(18) <= (i_crc(4) xor i_crc(5) xor i_crc(7) xor i_crc(26) xor i_data(4) xor i_data(5) xor i_data(7));
  s_result8(19) <= (i_crc(0) xor i_crc(1) xor i_crc(2) xor i_crc(3) xor i_crc(4) xor i_crc(5) xor i_crc(6) xor i_crc(27) xor i_data(0) xor i_data(1) xor i_data(2) xor i_data(3) xor i_data(4) xor i_data(5) xor i_data(6));
  s_result8(20) <= (i_crc(1) xor i_crc(2) xor i_crc(3) xor i_crc(4) xor i_crc(5) xor i_crc(6) xor i_crc(7) xor i_crc(28) xor i_data(1) xor i_data(2) xor i_data(3) xor i_data(4) xor i_data(5) xor i_data(6) xor i_data(7));
  s_result8(21) <= (i_crc(0) xor i_crc(1) xor i_crc(5) xor i_crc(6) xor i_crc(7) xor i_crc(29) xor i_data(0) xor i_data(1) xor i_data(5) xor i_data(6) xor i_data(7));
  s_result8(22) <= (i_crc(0) xor i_crc(3) xor i_crc(4) xor i_crc(6) xor i_crc(7) xor i_crc(30) xor i_data(0) xor i_data(3) xor i_data(4) xor i_data(6) xor i_data(7));
  s_result8(23) <= (i_crc(2) xor i_crc(3) xor i_crc(5) xor i_crc(7) xor i_crc(31) xor i_data(2) xor i_data(3) xor i_data(5) xor i_data(7));
  s_result8(24) <= (i_crc(1) xor i_crc(2) xor i_crc(6) xor i_data(1) xor i_data(2) xor i_data(6));
  s_result8(25) <= (i_crc(0) xor i_crc(2) xor i_crc(3) xor i_crc(7) xor i_data(0) xor i_data(2) xor i_data(3) xor i_data(7));
  s_result8(26) <= (i_crc(2) xor i_data(2));
  s_result8(27) <= (i_crc(3) xor i_data(3));
  s_result8(28) <= (i_crc(0) xor i_crc(4) xor i_data(0) xor i_data(4));
  s_result8(29) <= (i_crc(0) xor i_crc(1) xor i_crc(5) xor i_data(0) xor i_data(1) xor i_data(5));
  s_result8(30) <= (i_crc(0) xor i_crc(1) xor i_crc(2) xor i_crc(6) xor i_data(0) xor i_data(1) xor i_data(2) xor i_data(6));
  s_result8(31) <= (i_crc(0) xor i_crc(1) xor i_crc(2) xor i_crc(3) xor i_crc(7) xor i_data(0) xor i_data(1) xor i_data(2) xor i_data(3) xor i_data(7));

  -- 16 bits per clock (only bits 15 downto 0 are used from i_data).
  s_result16(0) <= (i_crc(0) xor i_crc(4) xor i_crc(7) xor i_crc(8) xor i_crc(9) xor i_crc(10) xor i_crc(11) xor i_crc(12) xor i_crc(16) xor i_data(0) xor i_data(4) xor i_data(7) xor i_data(8) xor i_data(9) xor i_data(10) xor i_data(11) xor i_data(12));
  s_result16(1) <= (i_crc(0) xor i_crc(1) xor i_crc(5) xor i_crc(8) xor i_crc(9) xor i_crc(10) xor i_crc(11) xor i_crc(12) xor i_crc(13) xor i_crc(17) xor i_data(0) xor i_data(1) xor i_data(5) xor i_data(8) xor i_data(9) xor i_data(10) xor i_data(11) xor i_data(12) xor i_data(13));
  s_result16(2) <= (i_crc(0) xor i_crc(1) xor i_crc(2) xor i_crc(6) xor i_crc(9) xor i_crc(10) xor i_crc(11) xor i_crc(12) xor i_crc(13) xor i_crc(14) xor i_crc(18) xor i_data(0) xor i_data(1) xor i_data(2) xor i_data(6) xor i_data(9) xor i_data(10) xor i_data(11) xor i_data(12) xor i_data(13) xor i_data(14));
  s_result16(3) <= (i_crc(1) xor i_crc(2) xor i_crc(3) xor i_crc(7) xor i_crc(10) xor i_crc(11) xor i_crc(12) xor i_crc(13) xor i_crc(14) xor i_crc(15) xor i_crc(19) xor i_data(1) xor i_data(2) xor i_data(3) xor i_data(7) xor i_data(10) xor i_data(11) xor i_data(12) xor i_data(13) xor i_data(14) xor i_data(15));
  s_result16(4) <= (i_crc(0) xor i_crc(2) xor i_crc(3) xor i_crc(7) xor i_crc(9) xor i_crc(10) xor i_crc(13) xor i_crc(14) xor i_crc(15) xor i_crc(20) xor i_data(0) xor i_data(2) xor i_data(3) xor i_data(7) xor i_data(9) xor i_data(10) xor i_data(13) xor i_data(14) xor i_data(15));
  s_result16(5) <= (i_crc(0) xor i_crc(1) xor i_crc(3) xor i_crc(7) xor i_crc(9) xor i_crc(12) xor i_crc(14) xor i_crc(15) xor i_crc(21) xor i_data(0) xor i_data(1) xor i_data(3) xor i_data(7) xor i_data(9) xor i_data(12) xor i_data(14) xor i_data(15));
  s_result16(6) <= (i_crc(0) xor i_crc(1) xor i_crc(2) xor i_crc(7) xor i_crc(9) xor i_crc(11) xor i_crc(12) xor i_crc(13) xor i_crc(15) xor i_crc(22) xor i_data(0) xor i_data(1) xor i_data(2) xor i_data(7) xor i_data(9) xor i_data(11) xor i_data(12) xor i_data(13) xor i_data(15));
  s_result16(7) <= (i_crc(1) xor i_crc(2) xor i_crc(3) xor i_crc(4) xor i_crc(7) xor i_crc(9) xor i_crc(11) xor i_crc(13) xor i_crc(14) xor i_crc(23) xor i_data(1) xor i_data(2) xor i_data(3) xor i_data(4) xor i_data(7) xor i_data(9) xor i_data(11) xor i_data(13) xor i_data(14));
  s_result16(8) <= (i_crc(2) xor i_crc(3) xor i_crc(4) xor i_crc(5) xor i_crc(8) xor i_crc(10) xor i_crc(12) xor i_crc(14) xor i_crc(15) xor i_crc(24) xor i_data(2) xor i_data(3) xor i_data(4) xor i_data(5) xor i_data(8) xor i_data(10) xor i_data(12) xor i_data(14) xor i_data(15));
  s_result16(9) <= (i_crc(3) xor i_crc(5) xor i_crc(6) xor i_crc(7) xor i_crc(8) xor i_crc(10) xor i_crc(12) xor i_crc(13) xor i_crc(15) xor i_crc(25) xor i_data(3) xor i_data(5) xor i_data(6) xor i_data(7) xor i_data(8) xor i_data(10) xor i_data(12) xor i_data(13) xor i_data(15));
  s_result16(10) <= (i_crc(6) xor i_crc(10) xor i_crc(12) xor i_crc(13) xor i_crc(14) xor i_crc(26) xor i_data(6) xor i_data(10) xor i_data(12) xor i_data(13) xor i_data(14));
  s_result16(11) <= (i_crc(0) xor i_crc(7) xor i_crc(11) xor i_crc(13) xor i_crc(14) xor i_crc(15) xor i_crc(27) xor i_data(0) xor i_data(7) xor i_data(11) xor i_data(13) xor i_data(14) xor i_data(15));
  s_result16(12) <= (i_crc(0) xor i_crc(1) xor i_crc(4) xor i_crc(7) xor i_crc(9) xor i_crc(10) xor i_crc(11) xor i_crc(14) xor i_crc(15) xor i_crc(28) xor i_data(0) xor i_data(1) xor i_data(4) xor i_data(7) xor i_data(9) xor i_data(10) xor i_data(11) xor i_data(14) xor i_data(15));
  s_result16(13) <= (i_crc(1) xor i_crc(2) xor i_crc(4) xor i_crc(5) xor i_crc(7) xor i_crc(9) xor i_crc(15) xor i_crc(29) xor i_data(1) xor i_data(2) xor i_data(4) xor i_data(5) xor i_data(7) xor i_data(9) xor i_data(15));
  s_result16(14) <= (i_crc(2) xor i_crc(3) xor i_crc(4) xor i_crc(5) xor i_crc(6) xor i_crc(7) xor i_crc(9) xor i_crc(11) xor i_crc(12) xor i_crc(30) xor i_data(2) xor i_data(3) xor i_data(4) xor i_data(5) xor i_data(6) xor i_data(7) xor i_data(9) xor i_data(11) xor i_data(12));
  s_result16(15) <= (i_crc(0) xor i_crc(3) xor i_crc(4) xor i_crc(5) xor i_crc(6) xor i_crc(7) xor i_crc(8) xor i_crc(10) xor i_crc(12) xor i_crc(13) xor i_crc(31) xor i_data(0) xor i_data(3) xor i_data(4) xor i_data(5) xor i_data(6) xor i_data(7) xor i_data(8) xor i_data(10) xor i_data(12) xor i_data(13));
  s_result16(16) <= (i_crc(1) xor i_crc(4) xor i_crc(5) xor i_crc(6) xor i_crc(7) xor i_crc(8) xor i_crc(9) xor i_crc(11) xor i_crc(13) xor i_crc(14) xor i_data(1) xor i_data(4) xor i_data(5) xor i_data(6) xor i_data(7) xor i_data(8) xor i_data(9) xor i_data(11) xor i_data(13) xor i_data(14));
  s_result16(17) <= (i_crc(0) xor i_crc(2) xor i_crc(5) xor i_crc(6) xor i_crc(7) xor i_crc(8) xor i_crc(9) xor i_crc(10) xor i_crc(12) xor i_crc(14) xor i_crc(15) xor i_data(0) xor i_data(2) xor i_data(5) xor i_data(6) xor i_data(7) xor i_data(8) xor i_data(9) xor i_data(10) xor i_data(12) xor i_data(14) xor i_data(15));
  s_result16(18) <= (i_crc(1) xor i_crc(3) xor i_crc(4) xor i_crc(6) xor i_crc(12) xor i_crc(13) xor i_crc(15) xor i_data(1) xor i_data(3) xor i_data(4) xor i_data(6) xor i_data(12) xor i_data(13) xor i_data(15));
  s_result16(19) <= (i_crc(2) xor i_crc(5) xor i_crc(8) xor i_crc(9) xor i_crc(10) xor i_crc(11) xor i_crc(12) xor i_crc(13) xor i_crc(14) xor i_data(2) xor i_data(5) xor i_data(8) xor i_data(9) xor i_data(10) xor i_data(11) xor i_data(12) xor i_data(13) xor i_data(14));
  s_result16(20) <= (i_crc(3) xor i_crc(6) xor i_crc(9) xor i_crc(10) xor i_crc(11) xor i_crc(12) xor i_crc(13) xor i_crc(14) xor i_crc(15) xor i_data(3) xor i_data(6) xor i_data(9) xor i_data(10) xor i_data(11) xor i_data(12) xor i_data(13) xor i_data(14) xor i_data(15));
  s_result16(21) <= (i_crc(0) xor i_crc(8) xor i_crc(9) xor i_crc(13) xor i_crc(14) xor i_crc(15) xor i_data(0) xor i_data(8) xor i_data(9) xor i_data(13) xor i_data(14) xor i_data(15));
  s_result16(22) <= (i_crc(1) xor i_crc(4) xor i_crc(7) xor i_crc(8) xor i_crc(11) xor i_crc(12) xor i_crc(14) xor i_crc(15) xor i_data(1) xor i_data(4) xor i_data(7) xor i_data(8) xor i_data(11) xor i_data(12) xor i_data(14) xor i_data(15));
  s_result16(23) <= (i_crc(0) xor i_crc(2) xor i_crc(4) xor i_crc(5) xor i_crc(7) xor i_crc(10) xor i_crc(11) xor i_crc(13) xor i_crc(15) xor i_data(0) xor i_data(2) xor i_data(4) xor i_data(5) xor i_data(7) xor i_data(10) xor i_data(11) xor i_data(13) xor i_data(15));
  s_result16(24) <= (i_crc(0) xor i_crc(1) xor i_crc(3) xor i_crc(4) xor i_crc(5) xor i_crc(6) xor i_crc(7) xor i_crc(9) xor i_crc(10) xor i_crc(14) xor i_data(0) xor i_data(1) xor i_data(3) xor i_data(4) xor i_data(5) xor i_data(6) xor i_data(7) xor i_data(9) xor i_data(10) xor i_data(14));
  s_result16(25) <= (i_crc(0) xor i_crc(1) xor i_crc(2) xor i_crc(4) xor i_crc(5) xor i_crc(6) xor i_crc(7) xor i_crc(8) xor i_crc(10) xor i_crc(11) xor i_crc(15) xor i_data(0) xor i_data(1) xor i_data(2) xor i_data(4) xor i_data(5) xor i_data(6) xor i_data(7) xor i_data(8) xor i_data(10) xor i_data(11) xor i_data(15));
  s_result16(26) <= (i_crc(1) xor i_crc(2) xor i_crc(3) xor i_crc(4) xor i_crc(5) xor i_crc(6) xor i_crc(10) xor i_data(1) xor i_data(2) xor i_data(3) xor i_data(4) xor i_data(5) xor i_data(6) xor i_data(10));
  s_result16(27) <= (i_crc(2) xor i_crc(3) xor i_crc(4) xor i_crc(5) xor i_crc(6) xor i_crc(7) xor i_crc(11) xor i_data(2) xor i_data(3) xor i_data(4) xor i_data(5) xor i_data(6) xor i_data(7) xor i_data(11));
  s_result16(28) <= (i_crc(0) xor i_crc(3) xor i_crc(4) xor i_crc(5) xor i_crc(6) xor i_crc(7) xor i_crc(8) xor i_crc(12) xor i_data(0) xor i_data(3) xor i_data(4) xor i_data(5) xor i_data(6) xor i_data(7) xor i_data(8) xor i_data(12));
  s_result16(29) <= (i_crc(1) xor i_crc(4) xor i_crc(5) xor i_crc(6) xor i_crc(7) xor i_crc(8) xor i_crc(9) xor i_crc(13) xor i_data(1) xor i_data(4) xor i_data(5) xor i_data(6) xor i_data(7) xor i_data(8) xor i_data(9) xor i_data(13));
  s_result16(30) <= (i_crc(2) xor i_crc(5) xor i_crc(6) xor i_crc(7) xor i_crc(8) xor i_crc(9) xor i_crc(10) xor i_crc(14) xor i_data(2) xor i_data(5) xor i_data(6) xor i_data(7) xor i_data(8) xor i_data(9) xor i_data(10) xor i_data(14));
  s_result16(31) <= (i_crc(3) xor i_crc(6) xor i_crc(7) xor i_crc(8) xor i_crc(9) xor i_crc(10) xor i_crc(11) xor i_crc(15) xor i_data(3) xor i_data(6) xor i_data(7) xor i_data(8) xor i_data(9) xor i_data(10) xor i_data(11) xor i_data(15));

  -- 32 bits per clock.
  s_result32(0) <= (i_crc(1) xor i_crc(2) xor i_crc(4) xor i_crc(5) xor i_crc(6) xor i_crc(7) xor i_crc(9) xor i_crc(11) xor i_crc(14) xor i_crc(15) xor i_crc(16) xor i_crc(20) xor i_crc(23) xor i_crc(24) xor i_crc(25) xor i_crc(26) xor i_crc(27) xor i_crc(28) xor i_data(1) xor i_data(2) xor i_data(4) xor i_data(5) xor i_data(6) xor i_data(7) xor i_data(9) xor i_data(11) xor i_data(14) xor i_data(15) xor i_data(16) xor i_data(20) xor i_data(23) xor i_data(24) xor i_data(25) xor i_data(26) xor i_data(27) xor i_data(28));
  s_result32(1) <= (i_crc(2) xor i_crc(3) xor i_crc(5) xor i_crc(6) xor i_crc(7) xor i_crc(8) xor i_crc(10) xor i_crc(12) xor i_crc(15) xor i_crc(16) xor i_crc(17) xor i_crc(21) xor i_crc(24) xor i_crc(25) xor i_crc(26) xor i_crc(27) xor i_crc(28) xor i_crc(29) xor i_data(2) xor i_data(3) xor i_data(5) xor i_data(6) xor i_data(7) xor i_data(8) xor i_data(10) xor i_data(12) xor i_data(15) xor i_data(16) xor i_data(17) xor i_data(21) xor i_data(24) xor i_data(25) xor i_data(26) xor i_data(27) xor i_data(28) xor i_data(29));
  s_result32(2) <= (i_crc(3) xor i_crc(4) xor i_crc(6) xor i_crc(7) xor i_crc(8) xor i_crc(9) xor i_crc(11) xor i_crc(13) xor i_crc(16) xor i_crc(17) xor i_crc(18) xor i_crc(22) xor i_crc(25) xor i_crc(26) xor i_crc(27) xor i_crc(28) xor i_crc(29) xor i_crc(30) xor i_data(3) xor i_data(4) xor i_data(6) xor i_data(7) xor i_data(8) xor i_data(9) xor i_data(11) xor i_data(13) xor i_data(16) xor i_data(17) xor i_data(18) xor i_data(22) xor i_data(25) xor i_data(26) xor i_data(27) xor i_data(28) xor i_data(29) xor i_data(30));
  s_result32(3) <= (i_crc(0) xor i_crc(4) xor i_crc(5) xor i_crc(7) xor i_crc(8) xor i_crc(9) xor i_crc(10) xor i_crc(12) xor i_crc(14) xor i_crc(17) xor i_crc(18) xor i_crc(19) xor i_crc(23) xor i_crc(26) xor i_crc(27) xor i_crc(28) xor i_crc(29) xor i_crc(30) xor i_crc(31) xor i_data(0) xor i_data(4) xor i_data(5) xor i_data(7) xor i_data(8) xor i_data(9) xor i_data(10) xor i_data(12) xor i_data(14) xor i_data(17) xor i_data(18) xor i_data(19) xor i_data(23) xor i_data(26) xor i_data(27) xor i_data(28) xor i_data(29) xor i_data(30) xor i_data(31));
  s_result32(4) <= (i_crc(0) xor i_crc(2) xor i_crc(4) xor i_crc(7) xor i_crc(8) xor i_crc(10) xor i_crc(13) xor i_crc(14) xor i_crc(16) xor i_crc(18) xor i_crc(19) xor i_crc(23) xor i_crc(25) xor i_crc(26) xor i_crc(29) xor i_crc(30) xor i_crc(31) xor i_data(0) xor i_data(2) xor i_data(4) xor i_data(7) xor i_data(8) xor i_data(10) xor i_data(13) xor i_data(14) xor i_data(16) xor i_data(18) xor i_data(19) xor i_data(23) xor i_data(25) xor i_data(26) xor i_data(29) xor i_data(30) xor i_data(31));
  s_result32(5) <= (i_crc(0) xor i_crc(2) xor i_crc(3) xor i_crc(4) xor i_crc(6) xor i_crc(7) xor i_crc(8) xor i_crc(16) xor i_crc(17) xor i_crc(19) xor i_crc(23) xor i_crc(25) xor i_crc(28) xor i_crc(30) xor i_crc(31) xor i_data(0) xor i_data(2) xor i_data(3) xor i_data(4) xor i_data(6) xor i_data(7) xor i_data(8) xor i_data(16) xor i_data(17) xor i_data(19) xor i_data(23) xor i_data(25) xor i_data(28) xor i_data(30) xor i_data(31));
  s_result32(6) <= (i_crc(2) xor i_crc(3) xor i_crc(6) xor i_crc(8) xor i_crc(11) xor i_crc(14) xor i_crc(15) xor i_crc(16) xor i_crc(17) xor i_crc(18) xor i_crc(23) xor i_crc(25) xor i_crc(27) xor i_crc(28) xor i_crc(29) xor i_crc(31) xor i_data(2) xor i_data(3) xor i_data(6) xor i_data(8) xor i_data(11) xor i_data(14) xor i_data(15) xor i_data(16) xor i_data(17) xor i_data(18) xor i_data(23) xor i_data(25) xor i_data(27) xor i_data(28) xor i_data(29) xor i_data(31));
  s_result32(7) <= (i_crc(0) xor i_crc(1) xor i_crc(2) xor i_crc(3) xor i_crc(5) xor i_crc(6) xor i_crc(11) xor i_crc(12) xor i_crc(14) xor i_crc(17) xor i_crc(18) xor i_crc(19) xor i_crc(20) xor i_crc(23) xor i_crc(25) xor i_crc(27) xor i_crc(29) xor i_crc(30) xor i_data(0) xor i_data(1) xor i_data(2) xor i_data(3) xor i_data(5) xor i_data(6) xor i_data(11) xor i_data(12) xor i_data(14) xor i_data(17) xor i_data(18) xor i_data(19) xor i_data(20) xor i_data(23) xor i_data(25) xor i_data(27) xor i_data(29) xor i_data(30));
  s_result32(8) <= (i_crc(1) xor i_crc(2) xor i_crc(3) xor i_crc(4) xor i_crc(6) xor i_crc(7) xor i_crc(12) xor i_crc(13) xor i_crc(15) xor i_crc(18) xor i_crc(19) xor i_crc(20) xor i_crc(21) xor i_crc(24) xor i_crc(26) xor i_crc(28) xor i_crc(30) xor i_crc(31) xor i_data(1) xor i_data(2) xor i_data(3) xor i_data(4) xor i_data(6) xor i_data(7) xor i_data(12) xor i_data(13) xor i_data(15) xor i_data(18) xor i_data(19) xor i_data(20) xor i_data(21) xor i_data(24) xor i_data(26) xor i_data(28) xor i_data(30) xor i_data(31));
  s_result32(9) <= (i_crc(0) xor i_crc(1) xor i_crc(3) xor i_crc(6) xor i_crc(8) xor i_crc(9) xor i_crc(11) xor i_crc(13) xor i_crc(15) xor i_crc(19) xor i_crc(21) xor i_crc(22) xor i_crc(23) xor i_crc(24) xor i_crc(26) xor i_crc(28) xor i_crc(29) xor i_crc(31) xor i_data(0) xor i_data(1) xor i_data(3) xor i_data(6) xor i_data(8) xor i_data(9) xor i_data(11) xor i_data(13) xor i_data(15) xor i_data(19) xor i_data(21) xor i_data(22) xor i_data(23) xor i_data(24) xor i_data(26) xor i_data(28) xor i_data(29) xor i_data(31));
  s_result32(10) <= (i_crc(5) xor i_crc(6) xor i_crc(10) xor i_crc(11) xor i_crc(12) xor i_crc(15) xor i_crc(22) xor i_crc(26) xor i_crc(28) xor i_crc(29) xor i_crc(30) xor i_data(5) xor i_data(6) xor i_data(10) xor i_data(11) xor i_data(12) xor i_data(15) xor i_data(22) xor i_data(26) xor i_data(28) xor i_data(29) xor i_data(30));
  s_result32(11) <= (i_crc(0) xor i_crc(6) xor i_crc(7) xor i_crc(11) xor i_crc(12) xor i_crc(13) xor i_crc(16) xor i_crc(23) xor i_crc(27) xor i_crc(29) xor i_crc(30) xor i_crc(31) xor i_data(0) xor i_data(6) xor i_data(7) xor i_data(11) xor i_data(12) xor i_data(13) xor i_data(16) xor i_data(23) xor i_data(27) xor i_data(29) xor i_data(30) xor i_data(31));
  s_result32(12) <= (i_crc(2) xor i_crc(4) xor i_crc(5) xor i_crc(6) xor i_crc(8) xor i_crc(9) xor i_crc(11) xor i_crc(12) xor i_crc(13) xor i_crc(15) xor i_crc(16) xor i_crc(17) xor i_crc(20) xor i_crc(23) xor i_crc(25) xor i_crc(26) xor i_crc(27) xor i_crc(30) xor i_crc(31) xor i_data(2) xor i_data(4) xor i_data(5) xor i_data(6) xor i_data(8) xor i_data(9) xor i_data(11) xor i_data(12) xor i_data(13) xor i_data(15) xor i_data(16) xor i_data(17) xor i_data(20) xor i_data(23) xor i_data(25) xor i_data(26) xor i_data(27) xor i_data(30) xor i_data(31));
  s_result32(13) <= (i_crc(0) xor i_crc(1) xor i_crc(2) xor i_crc(3) xor i_crc(4) xor i_crc(10) xor i_crc(11) xor i_crc(12) xor i_crc(13) xor i_crc(15) xor i_crc(17) xor i_crc(18) xor i_crc(20) xor i_crc(21) xor i_crc(23) xor i_crc(25) xor i_crc(31) xor i_data(0) xor i_data(1) xor i_data(2) xor i_data(3) xor i_data(4) xor i_data(10) xor i_data(11) xor i_data(12) xor i_data(13) xor i_data(15) xor i_data(17) xor i_data(18) xor i_data(20) xor i_data(21) xor i_data(23) xor i_data(25) xor i_data(31));
  s_result32(14) <= (i_crc(3) xor i_crc(6) xor i_crc(7) xor i_crc(9) xor i_crc(12) xor i_crc(13) xor i_crc(15) xor i_crc(18) xor i_crc(19) xor i_crc(20) xor i_crc(21) xor i_crc(22) xor i_crc(23) xor i_crc(25) xor i_crc(27) xor i_crc(28) xor i_data(3) xor i_data(6) xor i_data(7) xor i_data(9) xor i_data(12) xor i_data(13) xor i_data(15) xor i_data(18) xor i_data(19) xor i_data(20) xor i_data(21) xor i_data(22) xor i_data(23) xor i_data(25) xor i_data(27) xor i_data(28));
  s_result32(15) <= (i_crc(0) xor i_crc(4) xor i_crc(7) xor i_crc(8) xor i_crc(10) xor i_crc(13) xor i_crc(14) xor i_crc(16) xor i_crc(19) xor i_crc(20) xor i_crc(21) xor i_crc(22) xor i_crc(23) xor i_crc(24) xor i_crc(26) xor i_crc(28) xor i_crc(29) xor i_data(0) xor i_data(4) xor i_data(7) xor i_data(8) xor i_data(10) xor i_data(13) xor i_data(14) xor i_data(16) xor i_data(19) xor i_data(20) xor i_data(21) xor i_data(22) xor i_data(23) xor i_data(24) xor i_data(26) xor i_data(28) xor i_data(29));
  s_result32(16) <= (i_crc(0) xor i_crc(1) xor i_crc(5) xor i_crc(8) xor i_crc(9) xor i_crc(11) xor i_crc(14) xor i_crc(15) xor i_crc(17) xor i_crc(20) xor i_crc(21) xor i_crc(22) xor i_crc(23) xor i_crc(24) xor i_crc(25) xor i_crc(27) xor i_crc(29) xor i_crc(30) xor i_data(0) xor i_data(1) xor i_data(5) xor i_data(8) xor i_data(9) xor i_data(11) xor i_data(14) xor i_data(15) xor i_data(17) xor i_data(20) xor i_data(21) xor i_data(22) xor i_data(23) xor i_data(24) xor i_data(25) xor i_data(27) xor i_data(29) xor i_data(30));
  s_result32(17) <= (i_crc(1) xor i_crc(2) xor i_crc(6) xor i_crc(9) xor i_crc(10) xor i_crc(12) xor i_crc(15) xor i_crc(16) xor i_crc(18) xor i_crc(21) xor i_crc(22) xor i_crc(23) xor i_crc(24) xor i_crc(25) xor i_crc(26) xor i_crc(28) xor i_crc(30) xor i_crc(31) xor i_data(1) xor i_data(2) xor i_data(6) xor i_data(9) xor i_data(10) xor i_data(12) xor i_data(15) xor i_data(16) xor i_data(18) xor i_data(21) xor i_data(22) xor i_data(23) xor i_data(24) xor i_data(25) xor i_data(26) xor i_data(28) xor i_data(30) xor i_data(31));
  s_result32(18) <= (i_crc(0) xor i_crc(1) xor i_crc(3) xor i_crc(4) xor i_crc(5) xor i_crc(6) xor i_crc(9) xor i_crc(10) xor i_crc(13) xor i_crc(14) xor i_crc(15) xor i_crc(17) xor i_crc(19) xor i_crc(20) xor i_crc(22) xor i_crc(28) xor i_crc(29) xor i_crc(31) xor i_data(0) xor i_data(1) xor i_data(3) xor i_data(4) xor i_data(5) xor i_data(6) xor i_data(9) xor i_data(10) xor i_data(13) xor i_data(14) xor i_data(15) xor i_data(17) xor i_data(19) xor i_data(20) xor i_data(22) xor i_data(28) xor i_data(29) xor i_data(31));
  s_result32(19) <= (i_crc(9) xor i_crc(10) xor i_crc(18) xor i_crc(21) xor i_crc(24) xor i_crc(25) xor i_crc(26) xor i_crc(27) xor i_crc(28) xor i_crc(29) xor i_crc(30) xor i_data(9) xor i_data(10) xor i_data(18) xor i_data(21) xor i_data(24) xor i_data(25) xor i_data(26) xor i_data(27) xor i_data(28) xor i_data(29) xor i_data(30));
  s_result32(20) <= (i_crc(10) xor i_crc(11) xor i_crc(19) xor i_crc(22) xor i_crc(25) xor i_crc(26) xor i_crc(27) xor i_crc(28) xor i_crc(29) xor i_crc(30) xor i_crc(31) xor i_data(10) xor i_data(11) xor i_data(19) xor i_data(22) xor i_data(25) xor i_data(26) xor i_data(27) xor i_data(28) xor i_data(29) xor i_data(30) xor i_data(31));
  s_result32(21) <= (i_crc(1) xor i_crc(2) xor i_crc(4) xor i_crc(5) xor i_crc(6) xor i_crc(7) xor i_crc(9) xor i_crc(12) xor i_crc(14) xor i_crc(15) xor i_crc(16) xor i_crc(24) xor i_crc(25) xor i_crc(29) xor i_crc(30) xor i_crc(31) xor i_data(1) xor i_data(2) xor i_data(4) xor i_data(5) xor i_data(6) xor i_data(7) xor i_data(9) xor i_data(12) xor i_data(14) xor i_data(15) xor i_data(16) xor i_data(24) xor i_data(25) xor i_data(29) xor i_data(30) xor i_data(31));
  s_result32(22) <= (i_crc(0) xor i_crc(1) xor i_crc(3) xor i_crc(4) xor i_crc(8) xor i_crc(9) xor i_crc(10) xor i_crc(11) xor i_crc(13) xor i_crc(14) xor i_crc(17) xor i_crc(20) xor i_crc(23) xor i_crc(24) xor i_crc(27) xor i_crc(28) xor i_crc(30) xor i_crc(31) xor i_data(0) xor i_data(1) xor i_data(3) xor i_data(4) xor i_data(8) xor i_data(9) xor i_data(10) xor i_data(11) xor i_data(13) xor i_data(14) xor i_data(17) xor i_data(20) xor i_data(23) xor i_data(24) xor i_data(27) xor i_data(28) xor i_data(30) xor i_data(31));
  s_result32(23) <= (i_crc(6) xor i_crc(7) xor i_crc(10) xor i_crc(12) xor i_crc(16) xor i_crc(18) xor i_crc(20) xor i_crc(21) xor i_crc(23) xor i_crc(26) xor i_crc(27) xor i_crc(29) xor i_crc(31) xor i_data(6) xor i_data(7) xor i_data(10) xor i_data(12) xor i_data(16) xor i_data(18) xor i_data(20) xor i_data(21) xor i_data(23) xor i_data(26) xor i_data(27) xor i_data(29) xor i_data(31));
  s_result32(24) <= (i_crc(0) xor i_crc(1) xor i_crc(2) xor i_crc(4) xor i_crc(5) xor i_crc(6) xor i_crc(8) xor i_crc(9) xor i_crc(13) xor i_crc(14) xor i_crc(15) xor i_crc(16) xor i_crc(17) xor i_crc(19) xor i_crc(20) xor i_crc(21) xor i_crc(22) xor i_crc(23) xor i_crc(25) xor i_crc(26) xor i_crc(30) xor i_data(0) xor i_data(1) xor i_data(2) xor i_data(4) xor i_data(5) xor i_data(6) xor i_data(8) xor i_data(9) xor i_data(13) xor i_data(14) xor i_data(15) xor i_data(16) xor i_data(17) xor i_data(19) xor i_data(20) xor i_data(21) xor i_data(22) xor i_data(23) xor i_data(25) xor i_data(26) xor i_data(30));
  s_result32(25) <= (i_crc(1) xor i_crc(2) xor i_crc(3) xor i_crc(5) xor i_crc(6) xor i_crc(7) xor i_crc(9) xor i_crc(10) xor i_crc(14) xor i_crc(15) xor i_crc(16) xor i_crc(17) xor i_crc(18) xor i_crc(20) xor i_crc(21) xor i_crc(22) xor i_crc(23) xor i_crc(24) xor i_crc(26) xor i_crc(27) xor i_crc(31) xor i_data(1) xor i_data(2) xor i_data(3) xor i_data(5) xor i_data(6) xor i_data(7) xor i_data(9) xor i_data(10) xor i_data(14) xor i_data(15) xor i_data(16) xor i_data(17) xor i_data(18) xor i_data(20) xor i_data(21) xor i_data(22) xor i_data(23) xor i_data(24) xor i_data(26) xor i_data(27) xor i_data(31));
  s_result32(26) <= (i_crc(0) xor i_crc(1) xor i_crc(3) xor i_crc(5) xor i_crc(8) xor i_crc(9) xor i_crc(10) xor i_crc(14) xor i_crc(17) xor i_crc(18) xor i_crc(19) xor i_crc(20) xor i_crc(21) xor i_crc(22) xor i_crc(26) xor i_data(0) xor i_data(1) xor i_data(3) xor i_data(5) xor i_data(8) xor i_data(9) xor i_data(10) xor i_data(14) xor i_data(17) xor i_data(18) xor i_data(19) xor i_data(20) xor i_data(21) xor i_data(22) xor i_data(26));
  s_result32(27) <= (i_crc(0) xor i_crc(1) xor i_crc(2) xor i_crc(4) xor i_crc(6) xor i_crc(9) xor i_crc(10) xor i_crc(11) xor i_crc(15) xor i_crc(18) xor i_crc(19) xor i_crc(20) xor i_crc(21) xor i_crc(22) xor i_crc(23) xor i_crc(27) xor i_data(0) xor i_data(1) xor i_data(2) xor i_data(4) xor i_data(6) xor i_data(9) xor i_data(10) xor i_data(11) xor i_data(15) xor i_data(18) xor i_data(19) xor i_data(20) xor i_data(21) xor i_data(22) xor i_data(23) xor i_data(27));
  s_result32(28) <= (i_crc(0) xor i_crc(1) xor i_crc(2) xor i_crc(3) xor i_crc(5) xor i_crc(7) xor i_crc(10) xor i_crc(11) xor i_crc(12) xor i_crc(16) xor i_crc(19) xor i_crc(20) xor i_crc(21) xor i_crc(22) xor i_crc(23) xor i_crc(24) xor i_crc(28) xor i_data(0) xor i_data(1) xor i_data(2) xor i_data(3) xor i_data(5) xor i_data(7) xor i_data(10) xor i_data(11) xor i_data(12) xor i_data(16) xor i_data(19) xor i_data(20) xor i_data(21) xor i_data(22) xor i_data(23) xor i_data(24) xor i_data(28));
  s_result32(29) <= (i_crc(1) xor i_crc(2) xor i_crc(3) xor i_crc(4) xor i_crc(6) xor i_crc(8) xor i_crc(11) xor i_crc(12) xor i_crc(13) xor i_crc(17) xor i_crc(20) xor i_crc(21) xor i_crc(22) xor i_crc(23) xor i_crc(24) xor i_crc(25) xor i_crc(29) xor i_data(1) xor i_data(2) xor i_data(3) xor i_data(4) xor i_data(6) xor i_data(8) xor i_data(11) xor i_data(12) xor i_data(13) xor i_data(17) xor i_data(20) xor i_data(21) xor i_data(22) xor i_data(23) xor i_data(24) xor i_data(25) xor i_data(29));
  s_result32(30) <= (i_crc(0) xor i_crc(2) xor i_crc(3) xor i_crc(4) xor i_crc(5) xor i_crc(7) xor i_crc(9) xor i_crc(12) xor i_crc(13) xor i_crc(14) xor i_crc(18) xor i_crc(21) xor i_crc(22) xor i_crc(23) xor i_crc(24) xor i_crc(25) xor i_crc(26) xor i_crc(30) xor i_data(0) xor i_data(2) xor i_data(3) xor i_data(4) xor i_data(5) xor i_data(7) xor i_data(9) xor i_data(12) xor i_data(13) xor i_data(14) xor i_data(18) xor i_data(21) xor i_data(22) xor i_data(23) xor i_data(24) xor i_data(25) xor i_data(26) xor i_data(30));
  s_result32(31) <= (i_crc(0) xor i_crc(1) xor i_crc(3) xor i_crc(4) xor i_crc(5) xor i_crc(6) xor i_crc(8) xor i_crc(10) xor i_crc(13) xor i_crc(14) xor i_crc(15) xor i_crc(19) xor i_crc(22) xor i_crc(23) xor i_crc(24) xor i_crc(25) xor i_crc(26) xor i_crc(27) xor i_crc(31) xor i_data(0) xor i_data(1) xor i_data(3) xor i_data(4) xor i_data(5) xor i_data(6) xor i_data(8) xor i_data(10) xor i_data(13) xor i_data(14) xor i_data(15) xor i_data(19) xor i_data(22) xor i_data(23) xor i_data(24) xor i_data(25) xor i_data(26) xor i_data(27) xor i_data(31));

  TypeMux: with i_packed_mode select
    o_result <=
        s_result8  when "00",  -- crc32c.8
        s_result16 when "01",  -- crc32c.16
        s_result32 when "10",  -- crc32c.32
        (others => '-') when others;
end rtl;
